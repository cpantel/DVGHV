`timescale 1ns/1ps


/*
A clock divider in Verilog, using the cascading
flip-flop method.
*/

module clock_divider(
  input clk,
  input reset,
  output reg clk_div2,
  output reg clk_div4,
  output reg clk_div8,
  output reg clk_div16
);

  // simple ripple clock divider
  always @(posedge reset)
  begin
     clk_div2 <= 0;
     clk_div4 <= 0;
     clk_div8 <= 0;
     clk_div16 <= 0;
  end
  
  always @(posedge clk)
    clk_div2 <= ~clk_div2;

  always @(posedge clk_div2)
    clk_div4 <= ~clk_div4;

  always @(posedge clk_div4)
    clk_div8 <= ~clk_div8;

  always @(posedge clk_div8)
    clk_div16 <= ~clk_div16;

endmodule
